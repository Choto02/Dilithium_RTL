module verify (
    input [] pk,
    input [] rho,
    output 
);
    
    // fsm u_fsm (

    // );

    // SHA_core u_SHA_core (

    // );

    // NTT u_NTT (

    // );


endmodule